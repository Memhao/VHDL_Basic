ENTITY test_gates IS
END test_gates;


